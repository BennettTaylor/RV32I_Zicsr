`timescale 1ns / 1ps
`include "header.vh"

module csr(
    /* CSR module inputs */
    input wire i_clk, // CPU clock
    input wire i_rst_n // Active low reset

);

endmodule;
