`timescale 1ns / 1ps
`include "header.vh"

module forward(
    /* Forwarding unit inputs */
    input wire i_clk, // CPU clock
    input wire i_rst_n // Active low reset

);

endmodule;
