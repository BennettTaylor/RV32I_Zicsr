`timescale 1ns / 1ps
`include "header.vh"

module write_back(
    /* Write back stage inputs */
    input wire i_clk, // CPU clock
    input wire i_rst_n // Active low reset
);

endmodule;
