`timescale 1ns / 1ps
`include "header.vh"

module forward(
    // System Inputs
    input wire i_clk, // System clock
    input wire i_rst_n // Active low reset

);

endmodule;
